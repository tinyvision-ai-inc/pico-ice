module top (
  input ICE_2
);
endmodule
