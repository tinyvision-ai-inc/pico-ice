module top
